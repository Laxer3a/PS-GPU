// `define ULTRA
`define LAXER_STUFF
